//register offsets for the DUT
`define CSR 2'b00;
`define DPR 2'b01,
`define CMDR 2'b10,
`define FSMR 2'b11;