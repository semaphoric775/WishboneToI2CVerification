//fully implemented in later project

class i2cmb_coverage extends ncsu_component;

    function new(string name="");
        super.new(name);
    endfunction
endclass