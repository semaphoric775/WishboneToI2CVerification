class i2cmb_environment extends ncsu_object;
    `ncsu_register_object(i2cmb_environment)

    function new(string name="");
        super.new(name);
    endfunction
endclass