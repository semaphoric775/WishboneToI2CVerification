package types_pkg;

    typedef enum bit {WRITE=0, READ} i2c_op_t;

endpackage
