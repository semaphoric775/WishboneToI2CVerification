class i2cmb_coverage;
    //TODO
endclass