typedef enum bit {WRITE=0, READ} i2c_op_t;

