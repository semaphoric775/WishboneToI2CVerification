package i2cmb_env_pkg;
    `include "src/i2c_op_t.svh"
endpackage
