//fully implemented in later project

class i2cmb_coverage extends ncsu_object;
    `ncsu_register_object(i2cmb_coverage)

    function new(string name="");
        super.new(name);
    endfunction
endclass